// vgaClock.sv
// Convertido a SystemVerilog

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module vgaClock (
		input  logic  ref_clk_clk,        //      ref_clk.clk
		input  logic  ref_reset_reset,    //    ref_reset.reset
		output logic  reset_source_reset, // reset_source.reset
		output logic  vga_clk_clk         //      vga_clk.clk
	);

	vgaClock_video_pll_0 video_pll_0 (
		.ref_clk_clk        (ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (ref_reset_reset),    //    ref_reset.reset
		.vga_clk_clk        (vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (reset_source_reset)  // reset_source.reset
	);

endmodule