`include "../PC/pc.sv"
`include "../ALU/alu.sv"
`include "../REGISTER_UNIT/register_unit.sv"
